library verilog;
use verilog.vl_types.all;
entity cpu_vlg_check_tst is
    port(
        ALU_Input_1_out : in     vl_logic_vector(7 downto 0);
        ALU_Input_2_out : in     vl_logic_vector(7 downto 0);
        ALU_Result_out  : in     vl_logic_vector(7 downto 0);
        Branch_NE_out   : in     vl_logic;
        Branch_out      : in     vl_logic;
        EXMEM_ALU_Result_out: in     vl_logic_vector(7 downto 0);
        EXMEM_Register_Rd_out: in     vl_logic_vector(4 downto 0);
        EXMEM_RegWrite_out: in     vl_logic;
        ForwardA_out    : in     vl_logic_vector(1 downto 0);
        ForwardB_out    : in     vl_logic_vector(1 downto 0);
        HDU_MemWrite_out: in     vl_logic;
        HDU_RegWrite_out: in     vl_logic;
        IDEX_MemRead_out: in     vl_logic;
        IDEX_Register_Rs_out: in     vl_logic_vector(4 downto 0);
        IDEX_Register_Rt_out: in     vl_logic_vector(4 downto 0);
        IF_AddResult_out: in     vl_logic_vector(7 downto 0);
        IF_Branch_out   : in     vl_logic;
        IF_BranchNE_out : in     vl_logic;
        IF_Flush_out    : in     vl_logic;
        IF_PCPlus4_out  : in     vl_logic_vector(7 downto 0);
        IF_ReadData1_out: in     vl_logic_vector(7 downto 0);
        IF_ReadData2_out: in     vl_logic_vector(7 downto 0);
        IF_SignExtend_out: in     vl_logic_vector(7 downto 0);
        IF_Zero_out     : in     vl_logic_vector(7 downto 0);
        IFID_Register_Rs_out: in     vl_logic_vector(4 downto 0);
        IFID_Register_Rt_out: in     vl_logic_vector(4 downto 0);
        Instruction_out : in     vl_logic_vector(31 downto 0);
        Mem_Address_out : in     vl_logic_vector(7 downto 0);
        MemRead_out     : in     vl_logic;
        MemReadData_out : in     vl_logic_vector(7 downto 0);
        MEMWB_Read_Data_out: in     vl_logic_vector(7 downto 0);
        MEMWB_Register_Rd_out: in     vl_logic_vector(4 downto 0);
        MEMWB_RegWrite_out: in     vl_logic;
        MemWrite_Data_out: in     vl_logic_vector(7 downto 0);
        MemWrite_out    : in     vl_logic;
        PC              : in     vl_logic_vector(7 downto 0);
        Read_Data1_out  : in     vl_logic_vector(7 downto 0);
        Read_Data2_out  : in     vl_logic_vector(7 downto 0);
        RegWrite_out    : in     vl_logic;
        RegWriteData_out: in     vl_logic_vector(7 downto 0);
        STALL_out       : in     vl_logic;
        WriteRegister_out: in     vl_logic_vector(4 downto 0);
        Zero_out        : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end cpu_vlg_check_tst;
