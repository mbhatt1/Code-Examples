library verilog;
use verilog.vl_types.all;
entity cpu_vlg_vec_tst is
end cpu_vlg_vec_tst;
