library verilog;
use verilog.vl_types.all;
entity cpu is
    port(
        PC              : out    vl_logic_vector(7 downto 0);
        Instruction_out : out    vl_logic_vector(31 downto 0);
        Read_Data1_out  : out    vl_logic_vector(7 downto 0);
        Read_Data2_out  : out    vl_logic_vector(7 downto 0);
        ALU_Input_1_out : out    vl_logic_vector(7 downto 0);
        ALU_Input_2_out : out    vl_logic_vector(7 downto 0);
        ALU_Result_out  : out    vl_logic_vector(7 downto 0);
        Branch_out      : out    vl_logic;
        Branch_NE_out   : out    vl_logic;
        Zero_out        : out    vl_logic;
        MemRead_out     : out    vl_logic;
        MemReadData_out : out    vl_logic_vector(7 downto 0);
        MemWrite_out    : out    vl_logic;
        Mem_Address_out : out    vl_logic_vector(7 downto 0);
        MemWrite_Data_out: out    vl_logic_vector(7 downto 0);
        RegWrite_out    : out    vl_logic;
        WriteRegister_out: out    vl_logic_vector(4 downto 0);
        RegWriteData_out: out    vl_logic_vector(7 downto 0);
        EXMEM_RegWrite_out: out    vl_logic;
        EXMEM_ALU_Result_out: out    vl_logic_vector(7 downto 0);
        EXMEM_Register_Rd_out: out    vl_logic_vector(4 downto 0);
        MEMWB_RegWrite_out: out    vl_logic;
        MEMWB_Register_Rd_out: out    vl_logic_vector(4 downto 0);
        MEMWB_Read_Data_out: out    vl_logic_vector(7 downto 0);
        IDEX_Register_Rs_out: out    vl_logic_vector(4 downto 0);
        IDEX_Register_Rt_out: out    vl_logic_vector(4 downto 0);
        ForwardA_out    : out    vl_logic_vector(1 downto 0);
        ForwardB_out    : out    vl_logic_vector(1 downto 0);
        IDEX_MemRead_out: out    vl_logic;
        IFID_Register_Rs_out: out    vl_logic_vector(4 downto 0);
        IFID_Register_Rt_out: out    vl_logic_vector(4 downto 0);
        STALL_out       : out    vl_logic;
        HDU_RegWrite_out: out    vl_logic;
        HDU_MemWrite_out: out    vl_logic;
        IF_Flush_out    : out    vl_logic;
        IF_ReadData1_out: out    vl_logic_vector(7 downto 0);
        IF_ReadData2_out: out    vl_logic_vector(7 downto 0);
        IF_SignExtend_out: out    vl_logic_vector(7 downto 0);
        IF_Branch_out   : out    vl_logic;
        IF_BranchNE_out : out    vl_logic;
        IF_PCPlus4_out  : out    vl_logic_vector(7 downto 0);
        IF_AddResult_out: out    vl_logic_vector(7 downto 0);
        IF_Zero_out     : out    vl_logic_vector(7 downto 0);
        Clock           : in     vl_logic;
        Reset           : in     vl_logic
    );
end cpu;
